`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2019/12/23 18:35:31
// Design Name: 
// Module Name: parameter_package
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
/////////////////////////////////////////////////////////////////////////////////
package parameter_package;

parameter  DATA_WIDTH   = 8      ;              
parameter  K            = 3      ;              
parameter  ADDR_WIDTH   = 32     ;               
parameter  ROW_WIDTH    = 10     ;               
parameter  S            = 1      ; 
parameter  BATCH        = 2      ;     
parameter  PRECISION     = 4      ;
parameter  TEST_LAYER_COUNT =13    ;

//   conv_0 parameter  
//                               conv_layer://0   , 1     , 2    , 3   , 4    , 5 	, 6		, 7		, 8		, 9		, 10	, 11	, 12	, 13                        
parameter integer CONV_REAL_HOUT [0:13]   =  {224 , 224	, 224  , 112 , 112	, 56	, 56	, 56	, 28	, 28	, 28	, 14	, 14	, 14    };   
parameter integer CONV_REAL_HINT [0:13]   =  {224 , 224	, 224  , 112 , 112	, 56	, 56	, 56	, 28	, 28	, 28	, 14	, 14	, 14    };   
parameter integer CONV_C         [0:13]   =  {3   , 3	  , 64   , 64	 , 128	, 128	, 256	, 256	, 256	, 512	, 512	, 512	, 512	, 512   };   
parameter integer CONV_N         [0:13]   =  {3   , 64  , 64   , 128 , 128	, 256	, 256	, 256	, 512	, 512	, 512	, 512	, 512	, 512   };   
parameter integer CONV_Wh        [0:13]   =  {5   , 5	  , 1	   , 1	 , 2	  , 1	  , 2 	, 2	  , 1	  , 27	, 27	, 6	  , 6	  , 6     };   
parameter integer CONV_Ww        [0:13]   =  {4   , 4	  , 9	   , 29	 , 29	  , 29	, 29	, 29	, 29	, 15	, 15	, 17	, 17	, 17    };   
parameter integer CONV_Ih        [0:13]   =  {4   , 4	  , 9	   , 29	 , 29	  , 29	, 29	, 29	, 29	, 15	, 15	, 17	, 17	, 17    };   
parameter integer CONV_Iw        [0:13]   =  {1   , 1	  , 45   , 7	 , 7	  , 7	  , 7	  , 7	  , 7	  , 1	  , 1	  , 1	  , 1	  , 1     };   
parameter integer CONV_BI        [0:13]   =  {2   , 2   , 2    , 2   , 2	  , 2   , 2   , 2   , 2   , 2   , 2   , 2   , 2   , 2     };    
//Due to the time consuming of the transmission handshake, the recommended bi parameter is used to use 2 to improve transmission efficiency


/*
        conv_layer:// 1     , 2    , 3   , 4    , 5 	, 6		, 7		, 8		, 9		, 10	, 11	, 12	, 13    
 CONV_REAL_HOUT  =  [ 224	, 224  , 112 , 112	, 56	, 56	, 56	, 28	, 28	, 28	, 14	, 14	, 14    ];
 CONV_REAL_HINT  =  [ 224	, 224  , 112 , 112	, 56	, 56	, 56	, 28	, 28	, 28	, 14	, 14	, 14    ];            
 CONV_C          =  [ 3	    , 64   , 64	 , 128	, 128	, 256	, 256	, 256	, 512	, 512	, 512	, 512	, 512   ];
 CONV_N          =  [ 64    , 64   , 128 , 128	, 256	, 256	, 256	, 512	, 512	, 512	, 512	, 512	, 512   ];
 CONV_Wh         =  [ 5	    , 1	   , 1	 , 2	, 1	    , 2 	, 2	    , 1	    , 27	, 27	, 6	    , 6	    , 6     ];          
 CONV_Ww         =  [ 4	    , 9	   , 29	 , 29	, 29	, 29	, 29	, 29	, 15	, 15	, 17	, 17	, 17    ]; 
 CONV_Ih         =  [ 4	    , 9	   , 29	 , 29	, 29	, 29	, 29	, 29	, 15	, 15	, 17	, 17	, 17    ];
 CONV_Iw         =  [ 1	    , 45   , 7	 , 7	, 7	    , 7	    , 7	    , 7	    , 1	    , 1	    , 1	    , 1	    , 1     ];
 CONV_BI         =  [ 2     , 2    , 2   , 2	, 2     , 2     , 2     , 2     , 2     , 2     , 2     , 2     , 2     ]; 
 fm_in_1 = int8(25*(rand(CONV_REAL_HINT(1),CONV_REAL_HINT(1),CONV_C(1),BATCH)-0.5));
 weight_01 = int8(32*(rand(3,3,CONV_C(01),CONV_N(01))-0.5));
 weight_02 = int8(32*(rand(3,3,CONV_C(02),CONV_N(02))-0.5));
 weight_03 = int8(32*(rand(3,3,CONV_C(03),CONV_N(03))-0.5));
 weight_04 = int8(32*(rand(3,3,CONV_C(04),CONV_N(04))-0.5));
 weight_05 = int8(32*(rand(3,3,CONV_C(05),CONV_N(05))-0.5));
 weight_06 = int8(32*(rand(3,3,CONV_C(06),CONV_N(06))-0.5));
 weight_07 = int8(32*(rand(3,3,CONV_C(07),CONV_N(07))-0.5));
 weight_08 = int8(32*(rand(3,3,CONV_C(08),CONV_N(08))-0.5));
 weight_09 = int8(32*(rand(3,3,CONV_C(09),CONV_N(09))-0.5));
 weight_10 = int8(32*(rand(3,3,CONV_C(10),CONV_N(10))-0.5));
 weight_11 = int8(32*(rand(3,3,CONV_C(11),CONV_N(11))-0.5));
 weight_12 = int8(32*(rand(3,3,CONV_C(12),CONV_N(12))-0.5));
 weight_13 = int8(32*(rand(3,3,CONV_C(13),CONV_N(13))-0.5));
 
 [         fm_out_1,...
 fm_out_reshape_1_1,...
  weight_reshape2_1,...
   fm_in_reshape1_1]=conv_data_weight_generate(          fm_in_1,...
                                                          weight_01,...                                   
                                                  CONV_REAL_HINT (01),...                         
                                                          CONV_C (01),...                                 
                                                          CONV_N (01),...                                 
                                                         CONV_Wh (01),...                                
                                                         CONV_Ww (01),...                                
                                                         CONV_Ih (01),...                                
                                                         CONV_Iw (01),...                                
                                                           'conv_01_',...                                
                                                         BATCH);                                       
  [         fm_out_2,...                                                    
  fm_out_reshape_1_2,...                                                    
   weight_reshape2_2,...                                                    
    fm_in_reshape1_2]=conv_data_weight_generate(          fm_out_1,...       
                                                           weight_02,...    
                                                   CONV_REAL_HINT (02),...   
                                                           CONV_C (02),...   
                                                           CONV_N (02),...   
                                                          CONV_Wh (02),...   
                                                          CONV_Ww (02),...   
                                                          CONV_Ih (02),...   
                                                          CONV_Iw (02),...   
                                                            'conv_02_',...  
                                                          BATCH);           
  [fm_out_2_pool]=max_pooling(fm_out_2); 
   [         fm_out_3,...                                                  
   fm_out_reshape_1_3,...                                                  
    weight_reshape2_3,...                                                  
     fm_in_reshape1_3]=conv_data_weight_generate(          fm_out_2_pool,...    
                                                            weight_03,...  
                                                    CONV_REAL_HINT (03),... 
                                                            CONV_C (03),... 
                                                            CONV_N (03),... 
                                                           CONV_Wh (03),... 
                                                           CONV_Ww (03),... 
                                                           CONV_Ih (03),... 
                                                           CONV_Iw (03),... 
                                                             'conv_03_',...
                                                           BATCH);   
    [         fm_out_4,...                                                         
    fm_out_reshape_1_4,...                                                   
     weight_reshape2_4,...                                                   
      fm_in_reshape1_4]=conv_data_weight_generate(          fm_out_3,...
                                                             weight_04,...   
                                                     CONV_REAL_HINT (04),...  
                                                             CONV_C (04),...  
                                                             CONV_N (04),...  
                                                            CONV_Wh (04),...  
                                                            CONV_Ww (04),...  
                                                            CONV_Ih (04),...  
                                                            CONV_Iw (04),...  
                                                              'conv_04_',... 
                                                            BATCH);          
      
      [fm_out_4_pool]=max_pooling(fm_out_4);  
      [         fm_out_5,...                                                   
      fm_out_reshape_1_5,...                                                   
       weight_reshape2_5,...                                                   
        fm_in_reshape1_5]=conv_data_weight_generate(          fm_out_4_pool,...
                                                               weight_05,...   
                                                       CONV_REAL_HINT (05),...  
                                                               CONV_C (05),...  
                                                               CONV_N (05),...  
                                                              CONV_Wh (05),...  
                                                              CONV_Ww (05),...  
                                                              CONV_Ih (05),...  
                                                              CONV_Iw (05),...  
                                                                'conv_05_',... 
                                                              BATCH);  
      [         fm_out_6,...                                                                                                           
      fm_out_reshape_1_6,...                                                           
       weight_reshape2_6,...                                                   
        fm_in_reshape1_6]=conv_data_weight_generate(          fm_out_5,...
                                                               weight_06,...   
                                                       CONV_REAL_HINT (06),...  
                                                               CONV_C (06),...  
                                                               CONV_N (06),...  
                                                              CONV_Wh (06),...  
                                                              CONV_Ww (06),...  
                                                              CONV_Ih (06),...  
                                                              CONV_Iw (06),...  
                                                                'conv_06_',... 
                                                              BATCH); 
      [         fm_out_7,...                                                           
      fm_out_reshape_1_7,...                                                  
       weight_reshape2_7,...                                                  
        fm_in_reshape1_7]=conv_data_weight_generate(          fm_out_6,...    
                                                               weight_07,...  
                                                       CONV_REAL_HINT (07),... 
                                                               CONV_C (07),... 
                                                               CONV_N (07),... 
                                                              CONV_Wh (07),... 
                                                              CONV_Ww (07),... 
                                                              CONV_Ih (07),... 
                                                              CONV_Iw (07),... 
                                                                'conv_07_',...
                                                              BATCH);            
                                                              
                                                              
       [fm_out_7_pool]=max_pooling(fm_out_7);                                                       
       [         fm_out_8,...                                                                                                           
       fm_out_reshape_1_8,...                                                                                                           
        weight_reshape2_8,...                                                                                                           
         fm_in_reshape1_8]=conv_data_weight_generate(          fm_out_7_pool,...                                                             
                                                                 weight_08,...                                                           
                                                        CONV_REAL_HINT (08),...                                                         
                                                                CONV_C (08),...                                                         
                                                                CONV_N (08),...                                                         
                                                               CONV_Wh (08),...                                                         
                                                               CONV_Ww (08),...                                                         
                                                               CONV_Ih (08),...                                                         
                                                               CONV_Iw (08),...                                                         
                                                                  'conv_08_',...                                                         
                                                               BATCH);            
                                                               
        [         fm_out_9,...                                                                                                              
        fm_out_reshape_1_9,...                                                                                                              
         weight_reshape2_9,...                                                                                                              
          fm_in_reshape1_9]=conv_data_weight_generate(          fm_out_8,...                                                           
                                                                  weight_09,...                                                             
                                                         CONV_REAL_HINT (09),...                                                            
                                                                 CONV_C (09),...                                                            
                                                                 CONV_N (09),...                                                            
                                                                CONV_Wh (09),...                                                            
                                                                CONV_Ww (09),...                                                            
                                                                CONV_Ih (09),...                                                            
                                                                CONV_Iw (09),...                                                            
                                                                   'conv_09_',...                                                           
                                                                BATCH);                                                                     
                                                               
        [         fm_out_10,...                                                                                                                
        fm_out_reshape_1_10,...                                                                                                                
         weight_reshape2_10,...                                                                                                                
          fm_in_reshape1_10]=conv_data_weight_generate(          fm_out_9,...                                                             
                                                                  weight_10,...                                                               
                                                         CONV_REAL_HINT (10),...                                                              
                                                                 CONV_C (10),...                                                              
                                                                 CONV_N (10),...                                                              
                                                                CONV_Wh (10),...                                                              
                                                                CONV_Ww (10),...                                                                                                                    
                                                                CONV_Ih (10),...                                                             
                                                                CONV_Iw (10),...                                                             
                                                                   'conv_10_',...                                                            
                                                                BATCH);                                                                      
         
         [fm_out_10_pool]=max_pooling(fm_out_10);
         [         fm_out_11,...                                                      
         fm_out_reshape_1_11,...                                                      
          weight_reshape2_11,...                                                      
           fm_in_reshape1_11]=conv_data_weight_generate(          fm_out_10_pool,...   
                                                                   weight_11,...     
                                                          CONV_REAL_HINT (11),...    
                                                                  CONV_C (11),...    
                                                                  CONV_N (11),...    
                                                                 CONV_Wh (11),...    
                                                                 CONV_Ww (11),...    
                                                                 CONV_Ih (11),...    
                                                                 CONV_Iw (11),...    
                                                                    'conv_11_',...   
                                                                 BATCH);             
         
        
           [         fm_out_12,...                                                      
           fm_out_reshape_1_12,...                                                      
            weight_reshape2_12,...                                                      
             fm_in_reshape1_12]=conv_data_weight_generate(          fm_out_11,...  
                                                                     weight_12,...      
                                                            CONV_REAL_HINT (12),...     
                                                                    CONV_C (12),...     
                                                                    CONV_N (12),...     
                                                                   CONV_Wh (12),...     
                                                                   CONV_Ww (12),...     
                                                                   CONV_Ih (12),...     
                                                                   CONV_Iw (12),...     
                                                                      'conv_12_',...    
                                                                   BATCH);              
        
           [         fm_out_13,...                                                      
           fm_out_reshape_1_13,...                                                      
            weight_reshape2_13,...                                                      
             fm_in_reshape1_13]=conv_data_weight_generate(          fm_out_12,...  
                                                                     weight_13,...      
                                                            CONV_REAL_HINT (13),...     
                                                                    CONV_C (13),...     
                                                                    CONV_N (13),...     
                                                                   CONV_Wh (13),...     
                                                                   CONV_Ww (13),...     
                                                                   CONV_Ih (13),...     
                                                                   CONV_Iw (13),...     
                                                                      'conv_13_',...    
                                                                   BATCH);                                                                  
save('weight_fin.mat','fm_in_1',...
                       'weight_01',...
                       'weight_02',...
                       'weight_03',...
                       'weight_04',...
                       'weight_05',...
                       'weight_06',...
                       'weight_07',...
                       'weight_08',...
                       'weight_09',...
                       'weight_10',...
                       'weight_11',...
                       'weight_12',...
                       'weight_13');
//   conv_1 parameter        
parameter  CONV_1_REAL_HOUT    = 56    ;                
parameter  CONV_1_REAL_HINT    = 56    ;                
parameter  CONV_1_C            = 3      ;              
parameter  CONV_1_N            = 64     ;               
parameter  CONV_1_Wh           = 5      ;              
parameter  CONV_1_Ww           = 4      ;              
parameter  CONV_1_Ih           = 4      ;              
parameter  CONV_1_Iw           = 1      ;              
parameter  CONV_1_BI           = 2      ;    
//   conv_2 parameter        
parameter  CONV_2_REAL_HOUT    = 56    ;                
parameter  CONV_2_REAL_HINT    = 56    ;                
parameter  CONV_2_C            = 64     ;              
parameter  CONV_2_N            = 64     ;               
parameter  CONV_2_Wh           = 1      ;              
parameter  CONV_2_Ww           = 9      ;              
parameter  CONV_2_Ih           = 9      ;              
parameter  CONV_2_Iw           = 45     ;              
parameter  CONV_2_BI           = 2      ;    
//   conv_3 parameter POOLING        
parameter  CONV_3_REAL_HOUT    = 28    ;                
parameter  CONV_3_REAL_HINT    = 28    ;                
parameter  CONV_3_C            = 64     ;              
parameter  CONV_3_N            = 128    ;               
parameter  CONV_3_Wh           = 1      ;              
parameter  CONV_3_Ww           = 29     ;              
parameter  CONV_3_Ih           = 29     ;              
parameter  CONV_3_Iw           = 7      ;              
parameter  CONV_3_BI           = 2      ;    
//   conv_1 parameter        
parameter  CONV_1_REAL_HOUT    = 224    ;                
parameter  CONV_1_REAL_HINT    = 224    ;                
parameter  CONV_1_C            = 3      ;              
parameter  CONV_1_N            = 64     ;               
parameter  CONV_1_Wh           = 5      ;              
parameter  CONV_1_Ww           = 4      ;              
parameter  CONV_1_Ih           = 4      ;              
parameter  CONV_1_Iw           = 1      ;              
parameter  CONV_1_BI           = 2      ;    
//   conv_1 parameter        
parameter  CONV_1_REAL_HOUT    = 224    ;                
parameter  CONV_1_REAL_HINT    = 224    ;                
parameter  CONV_1_C            = 3      ;              
parameter  CONV_1_N            = 64     ;               
parameter  CONV_1_Wh           = 5      ;              
parameter  CONV_1_Ww           = 4      ;              
parameter  CONV_1_Ih           = 4      ;              
parameter  CONV_1_Iw           = 1      ;              
parameter  CONV_1_BI           = 2      ;    
//   conv_1 parameter        
parameter  CONV_1_REAL_HOUT    = 224    ;                
parameter  CONV_1_REAL_HINT    = 224    ;                
parameter  CONV_1_C            = 3      ;              
parameter  CONV_1_N            = 64     ;               
parameter  CONV_1_Wh           = 5      ;              
parameter  CONV_1_Ww           = 4      ;              
parameter  CONV_1_Ih           = 4      ;              
parameter  CONV_1_Iw           = 1      ;              
parameter  CONV_1_BI           = 2      ;    
 
 //   conv_1 parameter        
parameter  CONV_1_REAL_HOUT    = 224    ;                
parameter  CONV_1_REAL_HINT    = 224    ;                
parameter  CONV_1_C            = 3      ;              
parameter  CONV_1_N            = 64     ;               
parameter  CONV_1_Wh           = 5      ;              
parameter  CONV_1_Ww           = 4      ;              
parameter  CONV_1_Ih           = 4      ;              
parameter  CONV_1_Iw           = 1      ;              
parameter  CONV_1_BI           = 2      ;    
//   conv_1 parameter        
parameter  CONV_1_REAL_HOUT    = 224    ;                
parameter  CONV_1_REAL_HINT    = 224    ;                
parameter  CONV_1_C            = 3      ;              
parameter  CONV_1_N            = 64     ;               
parameter  CONV_1_Wh           = 5      ;              
parameter  CONV_1_Ww           = 4      ;              
parameter  CONV_1_Ih           = 4      ;              
parameter  CONV_1_Iw           = 1      ;              
parameter  CONV_1_BI           = 2      ;    
//   conv_1 parameter        
parameter  CONV_1_REAL_HOUT    = 224    ;                
parameter  CONV_1_REAL_HINT    = 224    ;                
parameter  CONV_1_C            = 3      ;              
parameter  CONV_1_N            = 64     ;               
parameter  CONV_1_Wh           = 5      ;              
parameter  CONV_1_Ww           = 4      ;              
parameter  CONV_1_Ih           = 4      ;              
parameter  CONV_1_Iw           = 1      ;              
parameter  CONV_1_BI           = 2      ;    
//   conv_1 parameter        
parameter  CONV_1_REAL_HOUT    = 224    ;                
parameter  CONV_1_REAL_HINT    = 224    ;                
parameter  CONV_1_C            = 3      ;              
parameter  CONV_1_N            = 64     ;               
parameter  CONV_1_Wh           = 5      ;              
parameter  CONV_1_Ww           = 4      ;              
parameter  CONV_1_Ih           = 4      ;              
parameter  CONV_1_Iw           = 1      ;              
parameter  CONV_1_BI           = 2      ;    
//   conv_1 parameter        
parameter  CONV_1_REAL_HOUT    = 224    ;                
parameter  CONV_1_REAL_HINT    = 224    ;                
parameter  CONV_1_C            = 3      ;              
parameter  CONV_1_N            = 64     ;               
parameter  CONV_1_Wh           = 5      ;              
parameter  CONV_1_Ww           = 4      ;              
parameter  CONV_1_Ih           = 4      ;              
parameter  CONV_1_Iw           = 1      ;              
parameter  CONV_1_BI           = 2      ;    
        
     */

endpackage